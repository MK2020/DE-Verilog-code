module mux32_two_to1(

ALU....